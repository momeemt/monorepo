package register_params;
  parameter int OPERAND_WIDTH = 32;
  parameter int REGISTER_DESCRIPTOR_WIDTH = 5;
  parameter int REGISTER_SIZE = 32;
endpackage
