module write_back (
    input logic clk,
    input logic rst,
    input logic valid_input,
    input logic stall_input
);

endmodule

